-------------------------------------------------------------------------------
-- Title      : tf wrapper
-- Project    : 
-------------------------------------------------------------------------------
-- File       : tf_wrapper.vhd
-- Author     : Michael Oshiro  <mco62@cornell.edu>
-- Company    : Cornell University
-- Created    : 2024-01-19
-- Last update: 2024-01-19
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: Simple module to pack/unpack SectorProcessor inputs into vectors
-------------------------------------------------------------------------------
-- Copyright (c) 2024 Cornell University
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2022-01-19  1.0      oshiro  Created
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

use work.memUtil_pkg.all;
use work.memUtil_aux_pkg.all;

entity tf_wrapper is
  port (
    clk                      : in  std_logic;
    reset                    : in  std_logic;
    IR_start                 : in  std_logic;
    IR_bx_in                 : in  std_logic_vector(2 downto 0);
    TP_bx_out_0              : out std_logic_vector(2 downto 0); 
    TP_bx_out_vld            : out std_logic;
    TP_done                  : out std_logic;
    DL_39_link_AV_dout       : in  t_arr_DL_39_DATA;
    DL_39_link_empty_neg     : in  t_arr_DL_39_1b;
    DL_39_link_read          : out t_arr_DL_39_1b
    );
end entity tf_wrapper;

architecture rtl of tf_wrapper is

begin  -- architecture rtl

  SectorProcessor_1 : entity work.SectorProcessor
    port map (
      clk                            => clk,
      reset                          => reset,
      IR_start                       => IR_start,
      IR_bx_in                       => IR_bx_in,
      TP_bx_out_0                    => TP_bx_out_0,
      TP_bx_out_vld                  => TP_bx_out_vld,
      TP_done                        => TP_done,
      DL_PS10G_1_A_link_AV_dout      => DL_39_link_AV_dout(PS10G_1_A),
      DL_PS10G_1_A_link_empty_neg    => DL_39_link_empty_neg(PS10G_1_A),
      DL_PS10G_1_A_link_read         => DL_39_link_read(PS10G_1_A),
      DL_PS10G_1_B_link_AV_dout      => DL_39_link_AV_dout(PS10G_1_B),
      DL_PS10G_1_B_link_empty_neg    => DL_39_link_empty_neg(PS10G_1_B),
      DL_PS10G_1_B_link_read         => DL_39_link_read(PS10G_1_B),
      DL_PS10G_2_A_link_AV_dout      => DL_39_link_AV_dout(PS10G_2_A),
      DL_PS10G_2_A_link_empty_neg    => DL_39_link_empty_neg(PS10G_2_A),
      DL_PS10G_2_A_link_read         => DL_39_link_read(PS10G_2_A),
      DL_PS10G_2_B_link_AV_dout      => DL_39_link_AV_dout(PS10G_2_B),
      DL_PS10G_2_B_link_empty_neg    => DL_39_link_empty_neg(PS10G_2_B),
      DL_PS10G_2_B_link_read         => DL_39_link_read(PS10G_2_B),
      DL_PS10G_3_A_link_AV_dout      => DL_39_link_AV_dout(PS10G_3_A),
      DL_PS10G_3_A_link_empty_neg    => DL_39_link_empty_neg(PS10G_3_A),
      DL_PS10G_3_A_link_read         => DL_39_link_read(PS10G_3_A),
      DL_PS10G_3_B_link_AV_dout      => DL_39_link_AV_dout(PS10G_3_B),
      DL_PS10G_3_B_link_empty_neg    => DL_39_link_empty_neg(PS10G_3_B),
      DL_PS10G_3_B_link_read         => DL_39_link_read(PS10G_3_B),
      DL_PS10G_4_A_link_AV_dout      => DL_39_link_AV_dout(PS10G_4_A),
      DL_PS10G_4_A_link_empty_neg    => DL_39_link_empty_neg(PS10G_4_A),
      DL_PS10G_4_A_link_read         => DL_39_link_read(PS10G_4_A),
      DL_PS10G_4_B_link_AV_dout      => DL_39_link_AV_dout(PS10G_4_B),
      DL_PS10G_4_B_link_empty_neg    => DL_39_link_empty_neg(PS10G_4_B),
      DL_PS10G_4_B_link_read         => DL_39_link_read(PS10G_4_B),
      DL_PS_1_A_link_AV_dout         => DL_39_link_AV_dout(PS_1_A),
      DL_PS_1_A_link_empty_neg       => DL_39_link_empty_neg(PS_1_A),
      DL_PS_1_A_link_read            => DL_39_link_read(PS_1_A),
      DL_PS_1_B_link_AV_dout         => DL_39_link_AV_dout(PS_1_B),
      DL_PS_1_B_link_empty_neg       => DL_39_link_empty_neg(PS_1_B),
      DL_PS_1_B_link_read            => DL_39_link_read(PS_1_B),
      DL_PS_2_A_link_AV_dout         => DL_39_link_AV_dout(PS_2_A),
      DL_PS_2_A_link_empty_neg       => DL_39_link_empty_neg(PS_2_A),
      DL_PS_2_A_link_read            => DL_39_link_read(PS_2_A),
      DL_PS_2_B_link_AV_dout         => DL_39_link_AV_dout(PS_2_B),
      DL_PS_2_B_link_empty_neg       => DL_39_link_empty_neg(PS_2_B),
      DL_PS_2_B_link_read            => DL_39_link_read(PS_2_B),
      DL_negPS10G_1_A_link_AV_dout   => DL_39_link_AV_dout(negPS10G_1_A),
      DL_negPS10G_1_A_link_empty_neg => DL_39_link_empty_neg(negPS10G_1_A),
      DL_negPS10G_1_A_link_read      => DL_39_link_read(negPS10G_1_A),
      DL_negPS10G_1_B_link_AV_dout   => DL_39_link_AV_dout(negPS10G_1_B),
      DL_negPS10G_1_B_link_empty_neg => DL_39_link_empty_neg(negPS10G_1_B),
      DL_negPS10G_1_B_link_read      => DL_39_link_read(negPS10G_1_B),
      DL_negPS10G_2_A_link_AV_dout   => DL_39_link_AV_dout(negPS10G_2_A),
      DL_negPS10G_2_A_link_empty_neg => DL_39_link_empty_neg(negPS10G_2_A),
      DL_negPS10G_2_A_link_read      => DL_39_link_read(negPS10G_2_A),
      DL_negPS10G_2_B_link_AV_dout   => DL_39_link_AV_dout(negPS10G_2_B),
      DL_negPS10G_2_B_link_empty_neg => DL_39_link_empty_neg(negPS10G_2_B),
      DL_negPS10G_2_B_link_read      => DL_39_link_read(negPS10G_2_B),
      DL_negPS10G_3_A_link_AV_dout   => DL_39_link_AV_dout(negPS10G_3_A),
      DL_negPS10G_3_A_link_empty_neg => DL_39_link_empty_neg(negPS10G_3_A),
      DL_negPS10G_3_A_link_read      => DL_39_link_read(negPS10G_3_A),
      DL_negPS10G_3_B_link_AV_dout   => DL_39_link_AV_dout(negPS10G_3_B),
      DL_negPS10G_3_B_link_empty_neg => DL_39_link_empty_neg(negPS10G_3_B),
      DL_negPS10G_3_B_link_read      => DL_39_link_read(negPS10G_3_B),
      DL_negPS10G_4_A_link_AV_dout   => DL_39_link_AV_dout(negPS10G_4_A),
      DL_negPS10G_4_A_link_empty_neg => DL_39_link_empty_neg(negPS10G_4_A),
      DL_negPS10G_4_A_link_read      => DL_39_link_read(negPS10G_4_A),
      DL_negPS10G_4_B_link_AV_dout   => DL_39_link_AV_dout(negPS10G_4_B),
      DL_negPS10G_4_B_link_empty_neg => DL_39_link_empty_neg(negPS10G_4_B),
      DL_negPS10G_4_B_link_read      => DL_39_link_read(negPS10G_4_B),
      DL_negPS_1_A_link_AV_dout      => DL_39_link_AV_dout(negPS_1_A),
      DL_negPS_1_A_link_empty_neg    => DL_39_link_empty_neg(negPS_1_A),
      DL_negPS_1_A_link_read         => DL_39_link_read(negPS_1_A),
      DL_negPS_1_B_link_AV_dout      => DL_39_link_AV_dout(negPS_1_B),
      DL_negPS_1_B_link_empty_neg    => DL_39_link_empty_neg(negPS_1_B),
      DL_negPS_1_B_link_read         => DL_39_link_read(negPS_1_B),
      DL_negPS_2_A_link_AV_dout      => DL_39_link_AV_dout(negPS_2_A),
      DL_negPS_2_A_link_empty_neg    => DL_39_link_empty_neg(negPS_2_A),
      DL_negPS_2_A_link_read         => DL_39_link_read(negPS_2_A),
      DL_negPS_2_B_link_AV_dout      => DL_39_link_AV_dout(negPS_2_B),
      DL_negPS_2_B_link_empty_neg    => DL_39_link_empty_neg(negPS_2_B),
      DL_negPS_2_B_link_read         => DL_39_link_read(negPS_2_B),
      DL_twoS_1_A_link_AV_dout       => DL_39_link_AV_dout(twoS_1_A),
      DL_twoS_1_A_link_empty_neg     => DL_39_link_empty_neg(twoS_1_A),
      DL_twoS_1_A_link_read          => DL_39_link_read(twoS_1_A),
      DL_twoS_1_B_link_AV_dout       => DL_39_link_AV_dout(twoS_1_B),
      DL_twoS_1_B_link_empty_neg     => DL_39_link_empty_neg(twoS_1_B),
      DL_twoS_1_B_link_read          => DL_39_link_read(twoS_1_B),
      DL_twoS_2_A_link_AV_dout       => DL_39_link_AV_dout(twoS_2_A),
      DL_twoS_2_A_link_empty_neg     => DL_39_link_empty_neg(twoS_2_A),
      DL_twoS_2_A_link_read          => DL_39_link_read(twoS_2_A),
      DL_twoS_2_B_link_AV_dout       => DL_39_link_AV_dout(twoS_2_B),
      DL_twoS_2_B_link_empty_neg     => DL_39_link_empty_neg(twoS_2_B),
      DL_twoS_2_B_link_read          => DL_39_link_read(twoS_2_B),
      DL_twoS_3_A_link_AV_dout       => DL_39_link_AV_dout(twoS_3_A),
      DL_twoS_3_A_link_empty_neg     => DL_39_link_empty_neg(twoS_3_A),
      DL_twoS_3_A_link_read          => DL_39_link_read(twoS_3_A),
      DL_twoS_3_B_link_AV_dout       => DL_39_link_AV_dout(twoS_3_B),
      DL_twoS_3_B_link_empty_neg     => DL_39_link_empty_neg(twoS_3_B),
      DL_twoS_3_B_link_read          => DL_39_link_read(twoS_3_B),
      DL_twoS_4_A_link_AV_dout       => DL_39_link_AV_dout(twoS_4_A),
      DL_twoS_4_A_link_empty_neg     => DL_39_link_empty_neg(twoS_4_A),
      DL_twoS_4_A_link_read          => DL_39_link_read(twoS_4_A),
      DL_twoS_4_B_link_AV_dout       => DL_39_link_AV_dout(twoS_4_B),
      DL_twoS_4_B_link_empty_neg     => DL_39_link_empty_neg(twoS_4_B),
      DL_twoS_4_B_link_read          => DL_39_link_read(twoS_4_B),
      DL_twoS_5_A_link_AV_dout       => DL_39_link_AV_dout(twoS_5_A),
      DL_twoS_5_A_link_empty_neg     => DL_39_link_empty_neg(twoS_5_A),
      DL_twoS_5_A_link_read          => DL_39_link_read(twoS_5_A),
      DL_twoS_5_B_link_AV_dout       => DL_39_link_AV_dout(twoS_5_B),
      DL_twoS_5_B_link_empty_neg     => DL_39_link_empty_neg(twoS_5_B),
      DL_twoS_5_B_link_read          => DL_39_link_read(twoS_5_B),
      DL_twoS_6_A_link_AV_dout       => DL_39_link_AV_dout(twoS_6_A),
      DL_twoS_6_A_link_empty_neg     => DL_39_link_empty_neg(twoS_6_A),
      DL_twoS_6_A_link_read          => DL_39_link_read(twoS_6_A),
      DL_twoS_6_B_link_AV_dout       => DL_39_link_AV_dout(twoS_6_B),
      DL_twoS_6_B_link_empty_neg     => DL_39_link_empty_neg(twoS_6_B),
      DL_twoS_6_B_link_read          => DL_39_link_read(twoS_6_B),
      DL_neg2S_1_A_link_AV_dout      => DL_39_link_AV_dout(neg2S_1_A),
      DL_neg2S_1_A_link_empty_neg    => DL_39_link_empty_neg(neg2S_1_A),
      DL_neg2S_1_A_link_read         => DL_39_link_read(neg2S_1_A),
      DL_neg2S_1_B_link_AV_dout      => DL_39_link_AV_dout(neg2S_1_B),
      DL_neg2S_1_B_link_empty_neg    => DL_39_link_empty_neg(neg2S_1_B),
      DL_neg2S_1_B_link_read         => DL_39_link_read(neg2S_1_B),
      DL_neg2S_2_A_link_AV_dout      => DL_39_link_AV_dout(neg2S_2_A),
      DL_neg2S_2_A_link_empty_neg    => DL_39_link_empty_neg(neg2S_2_A),
      DL_neg2S_2_A_link_read         => DL_39_link_read(neg2S_2_A),
      DL_neg2S_2_B_link_AV_dout      => DL_39_link_AV_dout(neg2S_2_B),
      DL_neg2S_2_B_link_empty_neg    => DL_39_link_empty_neg(neg2S_2_B),
      DL_neg2S_2_B_link_read         => DL_39_link_read(neg2S_2_B),
      DL_neg2S_3_A_link_AV_dout      => DL_39_link_AV_dout(neg2S_3_A),
      DL_neg2S_3_A_link_empty_neg    => DL_39_link_empty_neg(neg2S_3_A),
      DL_neg2S_3_A_link_read         => DL_39_link_read(neg2S_3_A),
      DL_neg2S_3_B_link_AV_dout      => DL_39_link_AV_dout(neg2S_3_B),
      DL_neg2S_3_B_link_empty_neg    => DL_39_link_empty_neg(neg2S_3_B),
      DL_neg2S_3_B_link_read         => DL_39_link_read(neg2S_3_B),
      DL_neg2S_4_A_link_AV_dout      => DL_39_link_AV_dout(neg2S_4_A),
      DL_neg2S_4_A_link_empty_neg    => DL_39_link_empty_neg(neg2S_4_A),
      DL_neg2S_4_A_link_read         => DL_39_link_read(neg2S_4_A),
      DL_neg2S_4_B_link_AV_dout      => DL_39_link_AV_dout(neg2S_4_B),
      DL_neg2S_4_B_link_empty_neg    => DL_39_link_empty_neg(neg2S_4_B),
      DL_neg2S_4_B_link_read         => DL_39_link_read(neg2S_4_B),
      DL_neg2S_5_A_link_AV_dout      => DL_39_link_AV_dout(neg2S_5_A),
      DL_neg2S_5_A_link_empty_neg    => DL_39_link_empty_neg(neg2S_5_A),
      DL_neg2S_5_A_link_read         => DL_39_link_read(neg2S_5_A),
      DL_neg2S_5_B_link_AV_dout      => DL_39_link_AV_dout(neg2S_5_B),
      DL_neg2S_5_B_link_empty_neg    => DL_39_link_empty_neg(neg2S_5_B),
      DL_neg2S_5_B_link_read         => DL_39_link_read(neg2S_5_B),
      DL_neg2S_6_A_link_AV_dout      => DL_39_link_AV_dout(neg2S_6_A),
      DL_neg2S_6_A_link_empty_neg    => DL_39_link_empty_neg(neg2S_6_A),
      DL_neg2S_6_A_link_read         => DL_39_link_read(neg2S_6_A),
      DL_neg2S_6_B_link_AV_dout      => DL_39_link_AV_dout(neg2S_6_B),
      DL_neg2S_6_B_link_empty_neg    => DL_39_link_empty_neg(neg2S_6_B),
      DL_neg2S_6_B_link_read         => DL_39_link_read(neg2S_6_B),
      AS_L1PHIAn1_enb          => '0',
      AS_L1PHIAn1_V_readaddr   => "0000000000",
      AS_L1PHIAn1_V_dout       => open,
      AS_L1PHIAn1_AV_dout_nent => open,
      AS_L1PHIBn1_enb          => '0',
      AS_L1PHIBn1_V_readaddr   => "0000000000",
      AS_L1PHIBn1_V_dout       => open,
      AS_L1PHIBn1_AV_dout_nent => open,
      AS_L1PHICn1_enb          => '0',
      AS_L1PHICn1_V_readaddr   => "0000000000",
      AS_L1PHICn1_V_dout       => open,
      AS_L1PHICn1_AV_dout_nent => open,
      AS_L1PHIDn1_enb          => '0',
      AS_L1PHIDn1_V_readaddr   => "0000000000",
      AS_L1PHIDn1_V_dout       => open,
      AS_L1PHIDn1_AV_dout_nent => open,
      AS_L1PHIEn1_enb          => '0',
      AS_L1PHIEn1_V_readaddr   => "0000000000",
      AS_L1PHIEn1_V_dout       => open,
      AS_L1PHIEn1_AV_dout_nent => open,
      AS_L1PHIFn1_enb          => '0',
      AS_L1PHIFn1_V_readaddr   => "0000000000",
      AS_L1PHIFn1_V_dout       => open,
      AS_L1PHIFn1_AV_dout_nent => open,
      AS_L1PHIGn1_enb          => '0',
      AS_L1PHIGn1_V_readaddr   => "0000000000",
      AS_L1PHIGn1_V_dout       => open,
      AS_L1PHIGn1_AV_dout_nent => open,
      AS_L1PHIHn1_enb          => '0',
      AS_L1PHIHn1_V_readaddr   => "0000000000",
      AS_L1PHIHn1_V_dout       => open,
      AS_L1PHIHn1_AV_dout_nent => open,
      AS_L2PHIAn1_enb          => '0',
      AS_L2PHIAn1_V_readaddr   => "0000000000",
      AS_L2PHIAn1_V_dout       => open,
      AS_L2PHIAn1_AV_dout_nent => open,
      AS_L2PHIBn1_enb          => '0',
      AS_L2PHIBn1_V_readaddr   => "0000000000",
      AS_L2PHIBn1_V_dout       => open,
      AS_L2PHIBn1_AV_dout_nent => open,
      AS_L2PHICn1_enb          => '0',
      AS_L2PHICn1_V_readaddr   => "0000000000",
      AS_L2PHICn1_V_dout       => open,
      AS_L2PHICn1_AV_dout_nent => open,
      AS_L2PHIDn1_enb          => '0',
      AS_L2PHIDn1_V_readaddr   => "0000000000",
      AS_L2PHIDn1_V_dout       => open,
      AS_L2PHIDn1_AV_dout_nent => open,
      AS_L3PHIAn1_enb          => '0',
      AS_L3PHIAn1_V_readaddr   => "0000000000",
      AS_L3PHIAn1_V_dout       => open,
      AS_L3PHIAn1_AV_dout_nent => open,
      AS_L3PHIBn1_enb          => '0',
      AS_L3PHIBn1_V_readaddr   => "0000000000",
      AS_L3PHIBn1_V_dout       => open,
      AS_L3PHIBn1_AV_dout_nent => open,
      AS_L3PHICn1_enb          => '0',
      AS_L3PHICn1_V_readaddr   => "0000000000",
      AS_L3PHICn1_V_dout       => open,
      AS_L3PHICn1_AV_dout_nent => open,
      AS_L3PHIDn1_enb          => '0',
      AS_L3PHIDn1_V_readaddr   => "0000000000",
      AS_L3PHIDn1_V_dout       => open,
      AS_L3PHIDn1_AV_dout_nent => open,
      AS_L4PHIAn1_enb          => '0',
      AS_L4PHIAn1_V_readaddr   => "0000000000",
      AS_L4PHIAn1_V_dout       => open,
      AS_L4PHIAn1_AV_dout_nent => open,
      AS_L4PHIBn1_enb          => '0',
      AS_L4PHIBn1_V_readaddr   => "0000000000",
      AS_L4PHIBn1_V_dout       => open,
      AS_L4PHIBn1_AV_dout_nent => open,
      AS_L4PHICn1_enb          => '0',
      AS_L4PHICn1_V_readaddr   => "0000000000",
      AS_L4PHICn1_V_dout       => open,
      AS_L4PHICn1_AV_dout_nent => open,
      AS_L4PHIDn1_enb          => '0',
      AS_L4PHIDn1_V_readaddr   => "0000000000",
      AS_L4PHIDn1_V_dout       => open,
      AS_L4PHIDn1_AV_dout_nent => open,
      AS_L5PHIAn1_enb          => '0',
      AS_L5PHIAn1_V_readaddr   => "0000000000",
      AS_L5PHIAn1_V_dout       => open,
      AS_L5PHIAn1_AV_dout_nent => open,
      AS_L5PHIBn1_enb          => '0',
      AS_L5PHIBn1_V_readaddr   => "0000000000",
      AS_L5PHIBn1_V_dout       => open,
      AS_L5PHIBn1_AV_dout_nent => open,
      AS_L5PHICn1_enb          => '0',
      AS_L5PHICn1_V_readaddr   => "0000000000",
      AS_L5PHICn1_V_dout       => open,
      AS_L5PHICn1_AV_dout_nent => open,
      AS_L5PHIDn1_enb          => '0',
      AS_L5PHIDn1_V_readaddr   => "0000000000",
      AS_L5PHIDn1_V_dout       => open,
      AS_L5PHIDn1_AV_dout_nent => open,
      AS_L6PHIAn1_enb          => '0',
      AS_L6PHIAn1_V_readaddr   => "0000000000",
      AS_L6PHIAn1_V_dout       => open,
      AS_L6PHIAn1_AV_dout_nent => open,
      AS_L6PHIBn1_enb          => '0',
      AS_L6PHIBn1_V_readaddr   => "0000000000",
      AS_L6PHIBn1_V_dout       => open,
      AS_L6PHIBn1_AV_dout_nent => open,
      AS_L6PHICn1_enb          => '0',
      AS_L6PHICn1_V_readaddr   => "0000000000",
      AS_L6PHICn1_V_dout       => open,
      AS_L6PHICn1_AV_dout_nent => open,
      AS_L6PHIDn1_enb          => '0',
      AS_L6PHIDn1_V_readaddr   => "0000000000",
      AS_L6PHIDn1_V_dout       => open,
      AS_L6PHIDn1_AV_dout_nent => open,
      AS_D1PHIAn1_enb          => '0',
      AS_D1PHIAn1_V_readaddr   => "0000000000",
      AS_D1PHIAn1_V_dout       => open,
      AS_D1PHIAn1_AV_dout_nent => open,
      AS_D1PHIBn1_enb          => '0',
      AS_D1PHIBn1_V_readaddr   => "0000000000",
      AS_D1PHIBn1_V_dout       => open,
      AS_D1PHIBn1_AV_dout_nent => open,
      AS_D1PHICn1_enb          => '0',
      AS_D1PHICn1_V_readaddr   => "0000000000",
      AS_D1PHICn1_V_dout       => open,
      AS_D1PHICn1_AV_dout_nent => open,
      AS_D1PHIDn1_enb          => '0',
      AS_D1PHIDn1_V_readaddr   => "0000000000",
      AS_D1PHIDn1_V_dout       => open,
      AS_D1PHIDn1_AV_dout_nent => open,
      AS_D2PHIAn1_enb          => '0',
      AS_D2PHIAn1_V_readaddr   => "0000000000",
      AS_D2PHIAn1_V_dout       => open,
      AS_D2PHIAn1_AV_dout_nent => open,
      AS_D2PHIBn1_enb          => '0',
      AS_D2PHIBn1_V_readaddr   => "0000000000",
      AS_D2PHIBn1_V_dout       => open,
      AS_D2PHIBn1_AV_dout_nent => open,
      AS_D2PHICn1_enb          => '0',
      AS_D2PHICn1_V_readaddr   => "0000000000",
      AS_D2PHICn1_V_dout       => open,
      AS_D2PHICn1_AV_dout_nent => open,
      AS_D2PHIDn1_enb          => '0',
      AS_D2PHIDn1_V_readaddr   => "0000000000",
      AS_D2PHIDn1_V_dout       => open,
      AS_D2PHIDn1_AV_dout_nent => open,
      AS_D3PHIAn1_enb          => '0',
      AS_D3PHIAn1_V_readaddr   => "0000000000",
      AS_D3PHIAn1_V_dout       => open,
      AS_D3PHIAn1_AV_dout_nent => open,
      AS_D3PHIBn1_enb          => '0',
      AS_D3PHIBn1_V_readaddr   => "0000000000",
      AS_D3PHIBn1_V_dout       => open,
      AS_D3PHIBn1_AV_dout_nent => open,
      AS_D3PHICn1_enb          => '0',
      AS_D3PHICn1_V_readaddr   => "0000000000",
      AS_D3PHICn1_V_dout       => open,
      AS_D3PHICn1_AV_dout_nent => open,
      AS_D3PHIDn1_enb          => '0',
      AS_D3PHIDn1_V_readaddr   => "0000000000",
      AS_D3PHIDn1_V_dout       => open,
      AS_D3PHIDn1_AV_dout_nent => open,
      AS_D4PHIAn1_enb          => '0',
      AS_D4PHIAn1_V_readaddr   => "0000000000",
      AS_D4PHIAn1_V_dout       => open,
      AS_D4PHIAn1_AV_dout_nent => open,
      AS_D4PHIBn1_enb          => '0',
      AS_D4PHIBn1_V_readaddr   => "0000000000",
      AS_D4PHIBn1_V_dout       => open,
      AS_D4PHIBn1_AV_dout_nent => open,
      AS_D4PHICn1_enb          => '0',
      AS_D4PHICn1_V_readaddr   => "0000000000",
      AS_D4PHICn1_V_dout       => open,
      AS_D4PHICn1_AV_dout_nent => open,
      AS_D4PHIDn1_enb          => '0',
      AS_D4PHIDn1_V_readaddr   => "0000000000",
      AS_D4PHIDn1_V_dout       => open,
      AS_D4PHIDn1_AV_dout_nent => open,
      AS_D5PHIAn1_enb          => '0',
      AS_D5PHIAn1_V_readaddr   => "0000000000",
      AS_D5PHIAn1_V_dout       => open,
      AS_D5PHIAn1_AV_dout_nent => open,
      AS_D5PHIBn1_enb          => '0',
      AS_D5PHIBn1_V_readaddr   => "0000000000",
      AS_D5PHIBn1_V_dout       => open,
      AS_D5PHIBn1_AV_dout_nent => open,
      AS_D5PHICn1_enb          => '0',
      AS_D5PHICn1_V_readaddr   => "0000000000",
      AS_D5PHICn1_V_dout       => open,
      AS_D5PHICn1_AV_dout_nent => open,
      AS_D5PHIDn1_enb          => '0',
      AS_D5PHIDn1_V_readaddr   => "0000000000",
      AS_D5PHIDn1_V_dout       => open,
      AS_D5PHIDn1_AV_dout_nent => open,
      TPAR_L1L2A_enb          => '0',
      TPAR_L1L2A_V_readaddr   => "0000000000",
      TPAR_L1L2A_V_dout       => open,
      TPAR_L1L2A_AV_dout_nent => open,
      TPAR_L1L2B_enb          => '0',
      TPAR_L1L2B_V_readaddr   => "0000000000",
      TPAR_L1L2B_V_dout       => open,
      TPAR_L1L2B_AV_dout_nent => open,
      TPAR_L1L2C_enb          => '0',
      TPAR_L1L2C_V_readaddr   => "0000000000",
      TPAR_L1L2C_V_dout       => open,
      TPAR_L1L2C_AV_dout_nent => open,
      TPAR_L1L2D_enb          => '0',
      TPAR_L1L2D_V_readaddr   => "0000000000",
      TPAR_L1L2D_V_dout       => open,
      TPAR_L1L2D_AV_dout_nent => open,
      TPAR_L1L2E_enb          => '0',
      TPAR_L1L2E_V_readaddr   => "0000000000",
      TPAR_L1L2E_V_dout       => open,
      TPAR_L1L2E_AV_dout_nent => open,
      TPAR_L1L2F_enb          => '0',
      TPAR_L1L2F_V_readaddr   => "0000000000",
      TPAR_L1L2F_V_dout       => open,
      TPAR_L1L2F_AV_dout_nent => open,
      TPAR_L1L2G_enb          => '0',
      TPAR_L1L2G_V_readaddr   => "0000000000",
      TPAR_L1L2G_V_dout       => open,
      TPAR_L1L2G_AV_dout_nent => open,
      TPAR_L1L2H_enb          => '0',
      TPAR_L1L2H_V_readaddr   => "0000000000",
      TPAR_L1L2H_V_dout       => open,
      TPAR_L1L2H_AV_dout_nent => open,
      TPAR_L1L2I_enb          => '0',
      TPAR_L1L2I_V_readaddr   => "0000000000",
      TPAR_L1L2I_V_dout       => open,
      TPAR_L1L2I_AV_dout_nent => open,
      TPAR_L1L2J_enb          => '0',
      TPAR_L1L2J_V_readaddr   => "0000000000",
      TPAR_L1L2J_V_dout       => open,
      TPAR_L1L2J_AV_dout_nent => open,
      TPAR_L1L2K_enb          => '0',
      TPAR_L1L2K_V_readaddr   => "0000000000",
      TPAR_L1L2K_V_dout       => open,
      TPAR_L1L2K_AV_dout_nent => open,
      TPAR_L1L2L_enb          => '0',
      TPAR_L1L2L_V_readaddr   => "0000000000",
      TPAR_L1L2L_V_dout       => open,
      TPAR_L1L2L_AV_dout_nent => open,
      TPAR_L2L3A_enb          => '0',
      TPAR_L2L3A_V_readaddr   => "0000000000",
      TPAR_L2L3A_V_dout       => open,
      TPAR_L2L3A_AV_dout_nent => open,
      TPAR_L2L3B_enb          => '0',
      TPAR_L2L3B_V_readaddr   => "0000000000",
      TPAR_L2L3B_V_dout       => open,
      TPAR_L2L3B_AV_dout_nent => open,
      TPAR_L2L3C_enb          => '0',
      TPAR_L2L3C_V_readaddr   => "0000000000",
      TPAR_L2L3C_V_dout       => open,
      TPAR_L2L3C_AV_dout_nent => open,
      TPAR_L2L3D_enb          => '0',
      TPAR_L2L3D_V_readaddr   => "0000000000",
      TPAR_L2L3D_V_dout       => open,
      TPAR_L2L3D_AV_dout_nent => open,
      TPAR_L3L4A_enb          => '0',
      TPAR_L3L4A_V_readaddr   => "0000000000",
      TPAR_L3L4A_V_dout       => open,
      TPAR_L3L4A_AV_dout_nent => open,
      TPAR_L3L4B_enb          => '0',
      TPAR_L3L4B_V_readaddr   => "0000000000",
      TPAR_L3L4B_V_dout       => open,
      TPAR_L3L4B_AV_dout_nent => open,
      TPAR_L3L4C_enb          => '0',
      TPAR_L3L4C_V_readaddr   => "0000000000",
      TPAR_L3L4C_V_dout       => open,
      TPAR_L3L4C_AV_dout_nent => open,
      TPAR_L3L4D_enb          => '0',
      TPAR_L3L4D_V_readaddr   => "0000000000",
      TPAR_L3L4D_V_dout       => open,
      TPAR_L3L4D_AV_dout_nent => open,
      TPAR_L5L6A_enb          => '0',
      TPAR_L5L6A_V_readaddr   => "0000000000",
      TPAR_L5L6A_V_dout       => open,
      TPAR_L5L6A_AV_dout_nent => open,
      TPAR_L5L6B_enb          => '0',
      TPAR_L5L6B_V_readaddr   => "0000000000",
      TPAR_L5L6B_V_dout       => open,
      TPAR_L5L6B_AV_dout_nent => open,
      TPAR_L5L6C_enb          => '0',
      TPAR_L5L6C_V_readaddr   => "0000000000",
      TPAR_L5L6C_V_dout       => open,
      TPAR_L5L6C_AV_dout_nent => open,
      TPAR_L5L6D_enb          => '0',
      TPAR_L5L6D_V_readaddr   => "0000000000",
      TPAR_L5L6D_V_dout       => open,
      TPAR_L5L6D_AV_dout_nent => open,
      TPAR_D1D2A_enb          => '0',
      TPAR_D1D2A_V_readaddr   => "0000000000",
      TPAR_D1D2A_V_dout       => open,
      TPAR_D1D2A_AV_dout_nent => open,
      TPAR_D1D2B_enb          => '0',
      TPAR_D1D2B_V_readaddr   => "0000000000",
      TPAR_D1D2B_V_dout       => open,
      TPAR_D1D2B_AV_dout_nent => open,
      TPAR_D1D2C_enb          => '0',
      TPAR_D1D2C_V_readaddr   => "0000000000",
      TPAR_D1D2C_V_dout       => open,
      TPAR_D1D2C_AV_dout_nent => open,
      TPAR_D1D2D_enb          => '0',
      TPAR_D1D2D_V_readaddr   => "0000000000",
      TPAR_D1D2D_V_dout       => open,
      TPAR_D1D2D_AV_dout_nent => open,
      TPAR_D3D4A_enb          => '0',
      TPAR_D3D4A_V_readaddr   => "0000000000",
      TPAR_D3D4A_V_dout       => open,
      TPAR_D3D4A_AV_dout_nent => open,
      TPAR_D3D4B_enb          => '0',
      TPAR_D3D4B_V_readaddr   => "0000000000",
      TPAR_D3D4B_V_dout       => open,
      TPAR_D3D4B_AV_dout_nent => open,
      TPAR_D3D4C_enb          => '0',
      TPAR_D3D4C_V_readaddr   => "0000000000",
      TPAR_D3D4C_V_dout       => open,
      TPAR_D3D4C_AV_dout_nent => open,
      TPAR_D3D4D_enb          => '0',
      TPAR_D3D4D_V_readaddr   => "0000000000",
      TPAR_D3D4D_V_dout       => open,
      TPAR_D3D4D_AV_dout_nent => open,
      TPAR_L1D1A_enb          => '0',
      TPAR_L1D1A_V_readaddr   => "0000000000",
      TPAR_L1D1A_V_dout       => open,
      TPAR_L1D1A_AV_dout_nent => open,
      TPAR_L1D1B_enb          => '0',
      TPAR_L1D1B_V_readaddr   => "0000000000",
      TPAR_L1D1B_V_dout       => open,
      TPAR_L1D1B_AV_dout_nent => open,
      TPAR_L1D1C_enb          => '0',
      TPAR_L1D1C_V_readaddr   => "0000000000",
      TPAR_L1D1C_V_dout       => open,
      TPAR_L1D1C_AV_dout_nent => open,
      TPAR_L1D1D_enb          => '0',
      TPAR_L1D1D_V_readaddr   => "0000000000",
      TPAR_L1D1D_V_dout       => open,
      TPAR_L1D1D_AV_dout_nent => open,
      TPAR_L1D1E_enb          => '0',
      TPAR_L1D1E_V_readaddr   => "0000000000",
      TPAR_L1D1E_V_dout       => open,
      TPAR_L1D1E_AV_dout_nent => open,
      TPAR_L1D1F_enb          => '0',
      TPAR_L1D1F_V_readaddr   => "0000000000",
      TPAR_L1D1F_V_dout       => open,
      TPAR_L1D1F_AV_dout_nent => open,
      TPAR_L1D1G_enb          => '0',
      TPAR_L1D1G_V_readaddr   => "0000000000",
      TPAR_L1D1G_V_dout       => open,
      TPAR_L1D1G_AV_dout_nent => open,
      TPAR_L1D1H_enb          => '0',
      TPAR_L1D1H_V_readaddr   => "0000000000",
      TPAR_L1D1H_V_dout       => open,
      TPAR_L1D1H_AV_dout_nent => open,
      TPAR_L2D1A_enb          => '0',
      TPAR_L2D1A_V_readaddr   => "0000000000",
      TPAR_L2D1A_V_dout       => open,
      TPAR_L2D1A_AV_dout_nent => open,
      TPAR_L2D1B_enb          => '0',
      TPAR_L2D1B_V_readaddr   => "0000000000",
      TPAR_L2D1B_V_dout       => open,
      TPAR_L2D1B_AV_dout_nent => open,
      TPAR_L2D1C_enb          => '0',
      TPAR_L2D1C_V_readaddr   => "0000000000",
      TPAR_L2D1C_V_dout       => open,
      TPAR_L2D1C_AV_dout_nent => open,
      TPAR_L2D1D_enb          => '0',
      TPAR_L2D1D_V_readaddr   => "0000000000",
      TPAR_L2D1D_V_dout       => open,
      TPAR_L2D1D_AV_dout_nent => open
      );

end architecture rtl;
